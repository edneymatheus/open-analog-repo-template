* Testbench: Smoke Test (Inverter)
* Path: sim/tb/tb_smoke.spice
*
* Goal: prove that a fresh clone can run ngspice from the repo root
* and write results into sim/results/ (ignored by git).

.include "../../ip/common/my_inverter.spice"

* Generic Level-1 MOS models (technology-agnostic)
.model nmos nmos level=1
.model pmos pmos level=1

.param VDD_VAL=1.8

VDD  vdd 0 {VDD_VAL}
VIN  in  0 PULSE(0 {VDD_VAL} 1n 100p 100p 10n 20n)

XINV in out vdd 0 my_inverter
CLOAD out 0 10f

.tran 50p 40n

.control
  set filetype=ascii
  run

  * Simple functional checks
  meas tran vout_max MAX v(out)
  meas tran vout_min MIN v(out)

  echo "Measured v(out):"
  print vout_max vout_min

  if (vout_max > 0.9*VDD_VAL) && (vout_min < 0.1*VDD_VAL)
    echo "TEST PASS: Inverter is switching!"
  else
    echo "TEST FAIL: Output did not swing rail-to-rail."
  end

  write "../results/smoke_test.raw" v(in) v(out)
  quit
.endc

.end
