* IP Block: Generic Inverter (Hello World)

.model nmos NMOS (LEVEL=1 VTO=0.6 KP=200u LAMBDA=0.02)
.model pmos PMOS (LEVEL=1 VTO=-0.6 KP=80u  LAMBDA=0.02)

.subckt my_inverter in out vdd gnd
M1 out in vdd vdd pmos w=2u l=0.5u
M2 out in gnd gnd nmos w=1u l=0.5u
.ends my_inverter
