* IP Block: Generic Inverter (Hello World)
* path: ip/common/my_inverter.spice

.subckt my_inverter in out vdd gnd
    Generic Ngspice model (level 1)
    M1 out in vdd vdd pmos w=2u l=0.5u
    M2 out in gnd gnd nmos w=1u l=0.5u
.ends my_inverter